module lab8_part_two (n,I,c,e,Q2,Q1,Q0);

	